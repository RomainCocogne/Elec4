
entity compteur is
	generic (N:	natural :=3);
	port (
		raz,h:	bit;
		q:	out bit_vector (N-1 downto 0)
	);
end entity;

architecture structure of compteur is
component bit0 is
	port(
		nraz,h:	bit;
		q0,c1:	out bit
	);
end component;
component biti is
	port(
		nraz,h,ci:	bit;
		qi,cip1:	out bit
	);
end component;

	signal c:	bit_vector(N downto 1);
	signal nraz:	bit;

begin
	cell0: bit0 port map (nraz,h,q(0),c(1));
	boucle: for i in 1 to (Q'high-1) generate
		celli: biti port map (nraz,h,c(i),q(i),c(i+1));
	end generate;

	nraz <= not raz;
end architecture;